`ifndef __RISCV_SV
`define __RISCV_SV

`ifdef VERILATOR
`include "include/common.sv"
`include "include/temp_storage.sv"

`include "src/regs.sv"

`include "src/IF/fetch.sv"
`include "src/ID/decoder.sv"
`include "src/EX/execute.sv"
`include "src/MEM/memory.sv"
`include "src/WB/writeback.sv"
`endif

module riscv
    import common::*;
    import temp_storage::*;
(
    // cpu basics
    input logic clk,
    input logic rst,

    // bus signals
	output ibus_req_t ireq,
	input ibus_resp_t iresp,

    // for DiffTest
    output word_t pc,
    output word_t [31:0] regs,
    output bool reg_write_enable,
	output reg_addr reg_dest_addr,
	output word_t reg_write_data,
	output bool valid,
	output inst_t inst,
	output addr_t inst_pc
);

	regs regs_inst (
		.clk(reg_write_clk),
		.rst(rst),
		.reg_write_enable(reg_write_enable),
		.reg_dest_addr(reg_dest_addr),
		.reg_write_data(reg_write_data),
		.regs_value(regs)
	);

	if_id if_id_state, if_id_state_new;
	id_ex id_ex_state, id_ex_state_new;
	ex_mem ex_mem_state, ex_mem_state_new;
	mem_wb mem_wb_state, mem_wb_state_new;

	bool fetch_inst_awaiting;

	bool awaiting = fetch_inst_awaiting;
	bool reg_write_clk;

    fetch fetch_instance (
		.ireq(ireq),
		.iresp(iresp),
		.pc(pc),
		.clk(clk),
		.rst(rst),
		.if_id_state(if_id_state_new),
		.awaiting(fetch_inst_awaiting)
    );

    decoder decoder_instance (
		// .clk(!awaiting ? clk : 0),
		// .clk(clk),

		.if_id_state(if_id_state),
		.id_ex_state(id_ex_state_new),

		.regs_value(regs),
		.rst(rst),
		.clk(reg_write_clk)
    );

    execute execute_instance (
		// .clk(!awaiting ? clk : 0),
		.clk(clk),

        .id_ex_state(id_ex_state),
        .ex_mem_state(ex_mem_state_new)
    );

	memory memory_instance (
		// .clk(!awaiting ? clk : 0),
		.clk(clk),

		.ex_mem_state(ex_mem_state),
		.mem_wb_state(mem_wb_state_new)
	);

	bool raw_valid_signal;
	bool delayed_1_clock_valid_signal;

	writeback writeback_instance (
		// .clk(!awaiting ? clk : 0),
		.clk(clk),

		.mem_wb_state(mem_wb_state),
		.reg_write_enable(reg_write_enable),
		.reg_dest_addr(reg_dest_addr),
		.reg_write_data(reg_write_data),

		.valid(raw_valid_signal),
		.inst(inst),
		.inst_pc(inst_pc),
		.reg_write_clk(reg_write_clk)
	);

	always_ff @(posedge clk or posedge rst) begin
		if (rst) begin
			// drink a cup of java ( also try brew! )
			// take on springboot
			// don't forget your redhat
		end else begin
			if_id_state <= if_id_state_new;
			id_ex_state <= id_ex_state_new;
			ex_mem_state <= ex_mem_state_new;
			mem_wb_state <= mem_wb_state_new;

			delayed_1_clock_valid_signal <= raw_valid_signal;
		end
	end

	assign valid = delayed_1_clock_valid_signal;

endmodule


`endif